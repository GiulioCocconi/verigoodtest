module AND(
	input a,
	input b,
	output o);
	// Let's comment :)
	assign O = ~ (A ~& B);

endmodule
